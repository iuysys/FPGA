library verilog;
use verilog.vl_types.all;
entity SR04_vlg_vec_tst is
end SR04_vlg_vec_tst;
