library verilog;
use verilog.vl_types.all;
entity SDRAM_tb is
end SDRAM_tb;
