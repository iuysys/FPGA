library verilog;
use verilog.vl_types.all;
entity CLK_DIV_EVEN_vlg_check_tst is
    port(
        CLK_OUT         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CLK_DIV_EVEN_vlg_check_tst;
