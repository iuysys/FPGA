library verilog;
use verilog.vl_types.all;
entity key_scan_vlg_vec_tst is
end key_scan_vlg_vec_tst;
