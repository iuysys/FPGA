library verilog;
use verilog.vl_types.all;
entity CLK_DIV_EVEN_vlg_vec_tst is
end CLK_DIV_EVEN_vlg_vec_tst;
