library verilog;
use verilog.vl_types.all;
entity UART_SDRAM_UART_tb is
end UART_SDRAM_UART_tb;
