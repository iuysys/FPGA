library verilog;
use verilog.vl_types.all;
entity UART_Txd_tb is
end UART_Txd_tb;
