library verilog;
use verilog.vl_types.all;
entity cycloneii_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end cycloneii_routing_wire;
