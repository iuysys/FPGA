library verilog;
use verilog.vl_types.all;
entity sdram_model_plus is
    generic(
        addr_bits       : integer := 12;
        data_bits       : integer := 16;
        col_bits        : integer := 8;
        mem_sizes       : integer := 1048575;
        tAC             : real    := 6.500000;
        tHZ             : real    := 5.500000;
        tOH             : integer := 2;
        tMRD            : real    := 2.000000;
        tRAS            : real    := 48.000000;
        tRC             : real    := 70.000000;
        tRCD            : real    := 20.000000;
        tRP             : real    := 20.000000;
        tRRD            : real    := 14.000000;
        tWRa            : real    := 7.500000;
        tWRp            : real    := 0.000000;
        Mode_Reg_Set    : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        Auto_Refresh    : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        Row_Active      : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        Pre_Charge      : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        PreCharge_All   : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        Write           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        Write_Pre       : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        Read            : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        Read_Pre        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        Burst_Stop      : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        Nop             : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        Dsel            : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1)
    );
    port(
        Dq              : inout  vl_logic_vector;
        Addr            : in     vl_logic_vector;
        Ba              : in     vl_logic_vector(1 downto 0);
        Clk             : in     vl_logic;
        Cke             : in     vl_logic;
        Cs_n            : in     vl_logic;
        Ras_n           : in     vl_logic;
        Cas_n           : in     vl_logic;
        We_n            : in     vl_logic;
        Dqm             : in     vl_logic_vector(3 downto 0);
        Debug           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of addr_bits : constant is 1;
    attribute mti_svvh_generic_type of data_bits : constant is 1;
    attribute mti_svvh_generic_type of col_bits : constant is 1;
    attribute mti_svvh_generic_type of mem_sizes : constant is 1;
    attribute mti_svvh_generic_type of tAC : constant is 1;
    attribute mti_svvh_generic_type of tHZ : constant is 1;
    attribute mti_svvh_generic_type of tOH : constant is 1;
    attribute mti_svvh_generic_type of tMRD : constant is 1;
    attribute mti_svvh_generic_type of tRAS : constant is 1;
    attribute mti_svvh_generic_type of tRC : constant is 1;
    attribute mti_svvh_generic_type of tRCD : constant is 1;
    attribute mti_svvh_generic_type of tRP : constant is 1;
    attribute mti_svvh_generic_type of tRRD : constant is 1;
    attribute mti_svvh_generic_type of tWRa : constant is 1;
    attribute mti_svvh_generic_type of tWRp : constant is 1;
    attribute mti_svvh_generic_type of Mode_Reg_Set : constant is 1;
    attribute mti_svvh_generic_type of Auto_Refresh : constant is 1;
    attribute mti_svvh_generic_type of Row_Active : constant is 1;
    attribute mti_svvh_generic_type of Pre_Charge : constant is 1;
    attribute mti_svvh_generic_type of PreCharge_All : constant is 1;
    attribute mti_svvh_generic_type of Write : constant is 1;
    attribute mti_svvh_generic_type of Write_Pre : constant is 1;
    attribute mti_svvh_generic_type of Read : constant is 1;
    attribute mti_svvh_generic_type of Read_Pre : constant is 1;
    attribute mti_svvh_generic_type of Burst_Stop : constant is 1;
    attribute mti_svvh_generic_type of Nop : constant is 1;
    attribute mti_svvh_generic_type of Dsel : constant is 1;
end sdram_model_plus;
