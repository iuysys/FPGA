library verilog;
use verilog.vl_types.all;
entity FIFO_T_vlg_tst is
end FIFO_T_vlg_tst;
