library verilog;
use verilog.vl_types.all;
entity washing_machine_vlg_vec_tst is
end washing_machine_vlg_vec_tst;
