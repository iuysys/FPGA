library verilog;
use verilog.vl_types.all;
entity SMG_vlg_vec_tst is
end SMG_vlg_vec_tst;
