library verilog;
use verilog.vl_types.all;
entity SDRAM_TOP_tb is
end SDRAM_TOP_tb;
