library verilog;
use verilog.vl_types.all;
entity washing_state_machine_vlg_vec_tst is
end washing_state_machine_vlg_vec_tst;
