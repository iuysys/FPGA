library verilog;
use verilog.vl_types.all;
entity OV7670_SDRAM_VGA_tb is
end OV7670_SDRAM_VGA_tb;
