library verilog;
use verilog.vl_types.all;
entity key_mod_vlg_vec_tst is
end key_mod_vlg_vec_tst;
