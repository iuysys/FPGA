module SMG(
	//输入
	CLK,RST_N,DATA,
	//输出
	SEL,DUAN
	
);
//-----------------------------------------------
//--外部信号
//-----------------------------------------------
input 				CLK;			
input 				RST_N;
input		[15:0] 	DATA;			//输入数据

output 	[2:0] 	SEL;			//位选信号端口
output 	[7:0] 	DUAN;			//段选信号端口
//-----------------------------------------------
//--内部信号
//-----------------------------------------------
reg 	[2:0] 	SEL_CNT;			//位选计数器		
reg 	[7:0] 	DUAN;				//段选数据端口寄存器
reg 	[7:0] 	DUAN_n;			//段选端口的下一个数据
//-----------------------------------------------
//-- 位选计数
//-----------------------------------------------
always@(posedge CLK or negedge RST_N)
begin
	if(!RST_N)
	begin
		SEL_CNT <= 3'b0;
	end
	else if(SEL_CNT == 3)
	begin
		SEL_CNT <= 3'b0;
	end
	else
		SEL_CNT <= SEL_CNT + 1'b1;
	
end
//-----------------------------------------------
//-- 输出位选信号
//-----------------------------------------------
assign SEL = SEL_CNT ;

//-----------------------------------------------
//-- 取出各位数据
//-----------------------------------------------
always@(SEL_CNT or DATA)
begin
	case(SEL_CNT)
		0	:
			DUAN_n <= DATA / 1_000 ;
		1	:
			DUAN_n <= DATA % 1_000 / 100 ;
		2	:
			DUAN_n <= DATA % 100 / 10 ;
		3	:
			DUAN_n <= DATA % 10 ;
		default :
			DUAN_n <= 8'b0 ;
	endcase
end
//-----------------------------------------------
//-- 输出段选信号
//-----------------------------------------------
always@(DUAN_n)
begin
	case(DUAN_n)
		0 : DUAN <=8'b00111111;//0
		1 : DUAN <=8'b00000110;//1
		2 : DUAN <=8'b01011011;//2
		3 : DUAN <=8'b01001111;//3
		4 : DUAN <=8'b01100110;//4
		5 : DUAN <=8'b01101101;//5
		6 : DUAN <=8'b01111101;//6
		7 : DUAN <=8'b00000111;//7
		8 : DUAN <=8'b01111111;//8
		9 : DUAN <=8'b01101111;//9
		default : 
			DUAN <= 8'b11111001;//E.
	endcase
end

endmodule















